-- adder/subtractor