library verilog;
use verilog.vl_types.all;
entity is_zero_vlg_vec_tst is
end is_zero_vlg_vec_tst;
