library verilog;
use verilog.vl_types.all;
entity is_zero_vlg_check_tst is
    port(
        ISZERO          : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end is_zero_vlg_check_tst;
